import JZJCoreFTypes::MemoryMode_t;

import EndiannessFunctions::toBigEndian32;
import EndiannessFunctions::toLittleEndian32;
import EndiannessFunctions::toBigEndian16;
import EndiannessFunctions::toLittleEndian16;

import BitExtensionFunctions::*;//todo specify only needed members

module MemoryController//2.5 port memory: 1 read port for instruction fetching, 1 read/write port for data loads/stores
#(
	parameter INITIAL_MEM_CONTENTS = "initialRam.mem",
	parameter RAM_A_WIDTH = 12
)
(
	input logic clock, reset,
	
	//Memory Mode and Control
	input MemoryMode_t memoryMode,//NOP will not allow error flags to be set
	input logic [2:0] funct3,
	
	//Addressing
	input logic [31:0] rs1,
	input logic [31:0] immediateI,
	input logic [31:0] immediateS,
	
	//Memory Loads
	output logic [31:0] memoryOutput,//Will only update if memoryMode is LOAD
	
	//Memory Stores
	input logic [31:0] rs2,//Will only write if memoryMode is STORE; for half words and bytes the memoryMode must be STORE_PRELOAD for 1 cycle first, then STORE to actually write
	
	//Instruction Fetching
	input logic [31:0] instructionAddressToAccess,
	output logic [31:0] instruction,
	
	//Error Flags
	output logic memoryUnalignedAccess,
	output logic memoryBadFunct3,
	
	//CPU memory mapped ports
	//Note that reads and writes are written to the addresses in little endian format
	//then converted back to be output / vise-versa for inputs
	//This makes it so for reads rd[0] = portXMemoryAddress[24] = portXInput[0]
	//and for writes............rs2[0] = portXMemoryAddress[24] = portXOutput[0]
	//My recomendation is therefore that ports are accessed whole words at a time
	//but if you keep the little endian -> big endian format in mind you can write half words or bytes
	//Reads from the address read from the input, writes write to the output
	//Inputs: (byte-wise read)				address (starting byte)
	input logic [31:0] portAInput,//		FFFFFFE0
	input logic [31:0] portBInput,//		FFFFFFE4
	input logic [31:0] portCInput,//   	FFFFFFE8
	input logic [31:0] portDInput,//   	FFFFFFEC
	input logic [31:0] portEInput,//   	FFFFFFF0
	input logic [31:0] portFInput,//   	FFFFFFF4
	input logic [31:0] portGInput,//   	FFFFFFF8
	input logic [31:0] portHInput,//   	FFFFFFFC
	//Outputs: (byte-wise write)			address (starting byte)
	output logic [31:0] portAOutput,//	FFFFFFE0
	output logic [31:0] portBOutput,//	FFFFFFE4
	output logic [31:0] portCOutput,//	FFFFFFE8
	output logic [31:0] portDOutput,//	FFFFFFEC
	output logic [31:0] portEOutput,//	FFFFFFF0
	output logic [31:0] portFOutput,//	FFFFFFF4
	output logic [31:0] portGOutput,//	FFFFFFF8
	output logic [31:0] portHOutput//	FFFFFFFC
	//For tristate ports, an additional port's outputs can be designated as a direction register, which can be used by and external module to allow/disalow writing
	//If feedback is desired, then inputs should be connected to their respective output register
	//MAKE SURE INPUTS ARE SYNCHRONIZED IF THEY ARE FROM ANOTHER CLOCK DOMAIN
);
/* Primitives */
//Addressing
logic [1:0] offset;
logic [31:0] addressToAccess;

//Backend Connections
logic [29:0] backendAddress;
logic [31:0] backendDataOut;
logic [31:0] backendDataIn;
logic backendWriteEnable;
logic [29:0] backendInstructionAddress;
logic [31:0] instructionLittleEndian;

assign backendWriteEnable = memoryMode == STORE;
assign instruction = toBigEndian32(instructionLittleEndian);

/* Addressing Logic */

assign backendInstructionAddress = instructionAddressToAccess[31:2];//If the instruction offset is bad, the ProgramCounter will set its error flag so we don't worry about that here

always_comb
begin
	case (memoryMode)
		LOAD: addressToAccess = rs1 + immediateI;
		STORE_PRELOAD, STORE: addressToAccess = rs1 + immediateS;//STORE_PRELOAD loads data currently at the address of the read-modify-write sequence
		default: addressToAccess = 'x;//Invalid enum
	endcase
end

assign backendAddress = addressToAccess[31:2];
assign offset = addressToAccess[1:0];

/* Modules */
//Internal
//Should be nested module but Quartus Prime does not support them :(
MemoryControllerLOADProcessor memoryControllerLOADProcessor(.*);
MemoryControllerSTOREProcessor memoryControllerSTOREProcessor(.*);
MemoryControllerErrorDetector errorDetector(.*);

//External
MemoryBackend #(.INITIAL_MEM_CONTENTS(INITIAL_MEM_CONTENTS), .RAM_A_WIDTH(RAM_A_WIDTH)) memoryBackend(.*);

endmodule: MemoryController

/* Internal Modules */

//Should be nested but Quartus Prime does not support nested modules :(
module MemoryControllerLOADProcessor
(
	//Inputs and raw memory data
	input logic [2:0] funct3,
	input logic [1:0] offset,
	input logic [31:0] backendDataOut,
	
	//Output (what to write to rd)
	output logic [31:0] memoryOutput
);
//backendDataOut to memoryOutput (reading/loading)
always_comb//Assumes memoryMode is LOAD since memoryOutput will be ignored anyways if it RDInputChooser has not selected memory
begin
	unique case (funct3)
		3'b000: memoryOutput = signExtend8To32(getByteAtOffset(backendDataOut, offset));//lb
		3'b001: memoryOutput = signExtend16To32(toBigEndian16(getHalfwordAtOffset(backendDataOut, offset)));//lh
		3'b010: memoryOutput = toBigEndian32(backendDataOut);//lw
		3'b100: memoryOutput = zeroExtend8To32(getByteAtOffset(backendDataOut, offset));//lbu
		3'b101: memoryOutput = zeroExtend16To32(toBigEndian16(getHalfwordAtOffset(backendDataOut, offset)));//lhu
		default: memoryOutput = 'x;//Bad funct3 or not LOAD
	endcase
end

//Selection Functions

function automatic logic [7:0] getByteAtOffset(input [31:0] data, input [1:0] offset);
begin
	unique case (offset)
		2'b00: getByteAtOffset = data[31:24];
		2'b01: getByteAtOffset = data[23:16];
		2'b10: getByteAtOffset = data[15:8];
		2'b11: getByteAtOffset = data[7:0];
	endcase
end
endfunction

function automatic logic [15:0] getHalfwordAtOffset(input [31:0] data, input [1:0] offset);
begin
	unique case (offset)
		2'b00: getHalfwordAtOffset = data[31:16];
		2'b10: getHalfwordAtOffset = data[15:0];
		default: getHalfwordAtOffset = 'x;//Bad offset
	endcase
end
endfunction

endmodule: MemoryControllerLOADProcessor

//Should be nested but Quartus Prime does not support nested modules :(
module MemoryControllerSTOREProcessor
(
	//Inputs, new data, and old raw memory data at the address to write to
	input logic [2:0] funct3,
	input logic [1:0] offset,
	input logic [31:0] rs2,
	input logic [31:0] backendDataOut,//old data
	
	//Output (what to write to the memory address)
	output logic [31:0] backendDataIn
);

//rs2 + (possibly) backendDataOut to backendDataIn (writing/storing)
always_comb//Assumes memoryMode is STORE since backendDataIn will not be writen unless memoryMode == STORE (see backendWriteEnable)
begin//If funct3 is sb or sh, backendDataOut will have already been updated with the original contents of an address last posedge (STORE_PRELOAD), so we can use that here
	unique case (funct3)
		3'b000: backendDataIn = replaceByteAtOffset(backendDataOut, rs2[7:0], offset);//sb
		3'b001: backendDataIn = replaceHalfwordAtOffset(backendDataOut, toLittleEndian16(rs2[15:0]), offset);//sh
		3'b010: backendDataIn = toLittleEndian32(rs2);//sw
		default: backendDataIn = 'x;//Bad funct3 or not STORE
	endcase
end

//Replacement Functions

function automatic logic [31:0] replaceByteAtOffset(input [31:0] data, input [7:0] newData, input [1:0] offset);
begin
	unique case (offset)
		2'b00: replaceByteAtOffset = {newData[7:0], data[23:0]};
		2'b01: replaceByteAtOffset = {data[31:24], newData[7:0], data[15:0]};
		2'b10: replaceByteAtOffset = {data[31:16], newData[7:0], data[7:0]};
		2'b11: replaceByteAtOffset = {data[31:8], newData[7:0]};
	endcase
end
endfunction

function automatic logic [31:0] replaceHalfwordAtOffset(input [31:0] data, input [15:0] newData, input [1:0] offset);
begin
	unique case (offset)
		2'b00: replaceHalfwordAtOffset = {newData[15:0], data[15:0]};
		2'b10: replaceHalfwordAtOffset = {data[31:16], newData[15:0]};
		default: replaceHalfwordAtOffset = 'x;//Bad offset
	endcase
end
endfunction

endmodule: MemoryControllerSTOREProcessor

//Should be nested but Quartus Prime does not support nested modules :(
module MemoryControllerErrorDetector
(
	//Inputs
	input MemoryMode_t memoryMode,
	input logic [2:0] funct3,
	input logic [1:0] offset,
	
	//Error Flags
	output logic memoryUnalignedAccess,
	output logic memoryBadFunct3
);

//Unaligned Access Detection
always_comb
begin
	unique case (memoryMode)
		LOAD, STORE_PRELOAD, STORE:
		begin
			unique case (funct3)
				3'b000, 3'b100: memoryUnalignedAccess = 1'b0;//lb/lbu | sb/Bad funct3
				3'b001, 3'b101: memoryUnalignedAccess = (offset == 2'b01) || (offset == 2'b11);//lh/lhu | sh/Bad funct3
				3'b010: memoryUnalignedAccess = offset != 2'b00;//lw | sw
				default: memoryUnalignedAccess = 1'bx;//Bad funct3
			endcase
		end
		NOP: memoryUnalignedAccess = 1'b0;//Not executing an instruction
		default: memoryUnalignedAccess = 1'bx;//Something is not right; bad enum
	endcase
end

//Bad Funct3 Detection
always_comb
begin
	unique case (memoryMode)
		LOAD: memoryBadFunct3 = (funct3 == 3'b011) || (funct3 == 3'b110)|| (funct3 == 3'b111);//None of these funct3s exist
		STORE_PRELOAD, STORE: memoryBadFunct3 = !((funct3 == 3'b000) || (funct3 == 3'b001)|| (funct3 == 3'b010));//Only these 3 funct3s exist
		NOP: memoryBadFunct3 = 1'b0;//Not executing an instruction
		default: memoryBadFunct3 = 1'bx;//Something is not right; bad enum
	endcase
end

endmodule: MemoryControllerErrorDetector