module MemoryBackend
(
	input clock, reset
	
	
);

endmodule 
